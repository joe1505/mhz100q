-- $Id: xilinx_2kx9_3e.vhd,v 1.2 2009/04/15 12:42:16 jrothwei Exp jrothwei $
-- Copyright 2009 Joseph Rothweiler
--------------------------------------------------------------------------------
-- Joseph Rothweiler, Sensicomm LLC, Branch 09Mar2009 from
-- d08_adcap/src/grabmem.vhd,v 1.1 2008/12/03 16:20:02
-- Using Xilinx Spartan 3E  internal block RAM as a 2k words x 9 bits RAM.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity xilinx_2kx9_3e is
    Port (
      clock1   : in  STD_LOGIC;
      write1   : in  STD_LOGIC;
      addr1    : in  STD_LOGIC_VECTOR (10 downto 0);
      data1in  : in  STD_LOGIC_VECTOR ( 8 downto 0);
      data1out : out STD_LOGIC_VECTOR ( 8 downto 0);
      --
      clock2   : in  STD_LOGIC;
      write2   : in  STD_LOGIC;
      addr2    : in  STD_LOGIC_VECTOR (10 downto 0);
      data2in  : in  STD_LOGIC_VECTOR ( 8 downto 0);
      data2out : out STD_LOGIC_VECTOR ( 8 downto 0)
    );
end xilinx_2kx9_3e;

architecture Behavioral of xilinx_2kx9_3e is
  signal CLKA  : std_logic;                     -- Port A Clock
  signal CLKB  : std_logic;                     -- Port B Clock
  signal DOA  : STD_LOGIC_VECTOR( 7 downto 0); -- A Data Output - lsb's used.
  signal DOB  : STD_LOGIC_VECTOR( 7 downto 0); -- B Data Output - lsb's used.
  signal DIA  : STD_LOGIC_VECTOR( 7 downto 0); -- A Data Input - lsb's used.
  signal DIB  : STD_LOGIC_VECTOR( 7 downto 0); -- B Data Input - lsb's used.
  signal DOPA : STD_LOGIC_VECTOR( 0 downto 0); -- A Parity Out. Unused.
  signal DOPB : STD_LOGIC_VECTOR( 0 downto 0); -- B Parity Out. Unused.
  signal DIPA : STD_LOGIC_VECTOR( 0 downto 0); -- A Parity In. Unused.
  signal DIPB : STD_LOGIC_VECTOR( 0 downto 0); -- B Parity In. Unused.
  signal ENA  : STD_LOGIC := '1';              -- A Enable. Not changed.
  signal ENB  : STD_LOGIC := '1';              -- B Enable. Not changed.
  signal SSRA : STD_LOGIC := '0';              -- A Sync Set/Reset. Not changed.
  signal SSRB : STD_LOGIC := '0';              -- B Sync Set/Reset. Not changed.
begin

   -- RAMB16_S9_S9: Virtex-II/II-Pro, Spartan-3/3E 2k x 8 + 1 Parity bit Dual-Port RAM
   -- Xilinx HDL Language Template, version 10.1.3


   RAMB16_S9_S9_inst : RAMB16_S9_S9
   generic map (
      INIT_A => X"000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Address 0 to 511
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 512 to 1023
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 1024 to 1535
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 1536 to 2047
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Address 0 to 511
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 512 to 1023
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 1024 to 1535
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 1536 to 2047
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
   )
   port map (
      DOA => DOA,      -- Port A 8-bit Data Output
      DOB => DOB,      -- Port B 8-bit Data Output
      DOPA => DOPA,    -- Port A 1-bit Parity Output
      DOPB => DOPB,    -- Port B 1-bit Parity Output
      ADDRA => addr1,  -- Port A 11-bit Address Input
      ADDRB => addr2,  -- Port B 11-bit Address Input
      CLKA => CLKA,    -- Port A Clock
      CLKB => CLKB,    -- Port B Clock
      DIA => DIA,      -- Port A 8-bit Data Input
      DIB => DIB,      -- Port B 8-bit Data Input
      DIPA => DIPA,    -- Port A 1-bit parity Input
      DIPB => DIPB,    -- Port-B 1-bit parity Input
      ENA => ENA,      -- Port A RAM Enable Input
      ENB => ENB,      -- PortB RAM Enable Input
      SSRA => SSRA,    -- Port A Synchronous Set/Reset Input
      SSRB => SSRB,    -- Port B Synchronous Set/Reset Input
      WEA => write1,   -- Port A Write Enable Input
      WEB => write2    -- Port B Write Enable Input
   );
   data1out <= DOPA & DOA;
   CLKA <= clock1;

   data2out <= DOPB & DOB;
   CLKB <= clock2;
   DIA <= data1in(7 downto 0);
   DIB <= data2in(7 downto 0);
   DIPA(0) <= data1in(8);
   DIPB(0) <= data2in(8);
end Behavioral;
